f<int> main() {
  printf("Hello World!");
}
